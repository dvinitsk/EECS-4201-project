// ----  Probes  ----
`define PROBE_ADDR      f_pc      //addr_i      
`define PROBE_DATA_IN   data_i    //mem_data_in
`define PROBE_DATA_OUT  data_o    //mem_data_out
`define PROBE_READ_EN   read_en   //mem_read_en
`define PROBE_WRITE_EN  write_en  //mem_write_en

`define PROBE_F_PC      f_pc    //fetch_pc_o
`define PROBE_F_INSN    f_inst  //fetch_insn_o 

// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
