// ----  Probes  ----
`define PROBE_ADDR      mem_addr
`define PROBE_DATA_IN   mem_data_in
`define PROBE_DATA_OUT  mem_data_out
`define PROBE_READ_EN   mem_read_en
`define PROBE_WRITE_EN  mem_write_en

`define PROBE_F_PC      fetch_pc_o
`define PROBE_F_INSN    fetch_insn_o //or change to mem_data_out 

// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd1
// ----  Top module  ----
